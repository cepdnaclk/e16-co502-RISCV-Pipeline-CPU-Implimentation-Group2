module ID_EX_pipeline_reg (
    ports
);


    
endmodule