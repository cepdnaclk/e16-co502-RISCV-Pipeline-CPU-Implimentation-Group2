`timescale  1ns/100ps
module ANDgate(IN1,IN2,OUT);
input IN1,IN2;
output OUT;
assign OUT = IN1 && IN2;
endmodule

